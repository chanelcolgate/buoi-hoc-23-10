parameter INTR_SFR_ADDR = 32'h400;
parameter CTRL_SFR_ADDR = 32'h404;
parameter IO_ADDR_SFR_ADDR = 32'h408;
parameter MEM_ADDR_SFR_ADDR = 32'h40C;
