class dpi_test extends test_base;
endclass
